// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
) (
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/

wire uart0_tx_wire;
wire uart1_tx_wire;

user_project mprj (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .wbs_sel_i(wbs_sel_i),
    .wbs_adr_i(wbs_adr_i),
    .wbs_dat_i(wbs_dat_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_dat_o(wbs_dat_o),
    .user_irq(user_irq),
    .uart0_rx(io_in[6]),
    .uart0_tx(uart0_tx_wire),
    .uart1_rx(io_in[8]),
    .uart1_tx(uart1_tx_wire)
);

assign io_out[0] = 1'b0;
assign io_oeb[0] = 1'b1;
assign io_out[1] = 1'b0;
assign io_oeb[1] = 1'b1;
assign io_out[2] = 1'b0;
assign io_oeb[2] = 1'b1;
assign io_out[3] = 1'b0;
assign io_oeb[3] = 1'b1;
assign io_out[4] = 1'b0;
assign io_oeb[4] = 1'b1;
assign io_out[5] = 1'b0;
assign io_oeb[5] = 1'b1;
assign io_out[6] = 1'b0;
assign io_oeb[6] = 1'b1;
assign io_out[7] = uart0_tx_wire;
assign io_oeb[7] = 1'b0;
assign io_out[8] = 1'b0;
assign io_oeb[8] = 1'b1;
assign io_out[9] = uart1_tx_wire;
assign io_oeb[9] = 1'b0;
assign io_out[10] = 1'b0;
assign io_oeb[10] = 1'b1;
assign io_out[11] = 1'b0;
assign io_oeb[11] = 1'b1;
assign io_out[12] = 1'b0;
assign io_oeb[12] = 1'b1;
assign io_out[13] = 1'b0;
assign io_oeb[13] = 1'b1;
assign io_out[14] = 1'b0;
assign io_oeb[14] = 1'b1;
assign io_out[15] = 1'b0;
assign io_oeb[15] = 1'b1;
assign io_out[16] = 1'b0;
assign io_oeb[16] = 1'b1;
assign io_out[17] = 1'b0;
assign io_oeb[17] = 1'b1;
assign io_out[18] = 1'b0;
assign io_oeb[18] = 1'b1;
assign io_out[19] = 1'b0;
assign io_oeb[19] = 1'b1;
assign io_out[20] = 1'b0;
assign io_oeb[20] = 1'b1;
assign io_out[21] = 1'b0;
assign io_oeb[21] = 1'b1;
assign io_out[22] = 1'b0;
assign io_oeb[22] = 1'b1;
assign io_out[23] = 1'b0;
assign io_oeb[23] = 1'b1;
assign io_out[24] = 1'b0;
assign io_oeb[24] = 1'b1;
assign io_out[25] = 1'b0;
assign io_oeb[25] = 1'b1;
assign io_out[26] = 1'b0;
assign io_oeb[26] = 1'b1;
assign io_out[27] = 1'b0;
assign io_oeb[27] = 1'b1;
assign io_out[28] = 1'b0;
assign io_oeb[28] = 1'b1;
assign io_out[29] = 1'b0;
assign io_oeb[29] = 1'b1;
assign io_out[30] = 1'b0;
assign io_oeb[30] = 1'b1;
assign io_out[31] = 1'b0;
assign io_oeb[31] = 1'b1;
assign io_out[32] = 1'b0;
assign io_oeb[32] = 1'b1;
assign io_out[33] = 1'b0;
assign io_oeb[33] = 1'b1;
assign io_out[34] = 1'b0;
assign io_oeb[34] = 1'b1;
assign io_out[35] = 1'b0;
assign io_oeb[35] = 1'b1;
assign io_out[36] = 1'b0;
assign io_oeb[36] = 1'b1;
assign io_out[37] = 1'b0;
assign io_oeb[37] = 1'b1;

assign la_data_out = 128'b0;

endmodule	// user_project_wrapper

`default_nettype wire
